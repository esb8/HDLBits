module top_module (
    input in1,
    input in2,
    output out
);
endmodule
